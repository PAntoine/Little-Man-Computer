--------------------------------------------------------------------------------
--                                                                 IO Controller
---                                                    LMC (Little Man Computer)
--------------------------------------------------------------------------------
--- Name:	io_controller.vhdl
--- Desc:
---       Little Man Computer
---	
---
--- Errors:
---       None.
---
--- Dependencies:
---       None.
---
--- Current Target: <don't know>
---
--- Author: Peter Antoine 
--- Date  : 17th Feb 2011
--------------------------------------------------------------------------------
---                                             Copyright (c) 2011 Peter Antoine
-----------------------------------------------------------------------------{{{
--- Version  Author  Date        Changes
--- -------  ------  ----------  ----------------------------------------------
--- 0.1      PA      17.02.2011  Initial Revision.
-----------------------------------------------------------------------------}}}


